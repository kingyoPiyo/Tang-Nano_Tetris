/********************************************************
* Title    : Character ROM
* Date     : 2019/10/22
* Design   : kingyo
********************************************************/
module char_rom (
    input   wire            i_clk,
    input   wire            i_res_n,
    input   wire    [ 5:0]  i_addr,
    output  reg     [63:0]  o_data
    )/* synthesis syn_romstyle = "block_rom" */;

    always @(posedge i_clk or negedge i_res_n) begin
        if (~i_res_n) begin
            o_data <= 64'd0;
        end else begin
            case (i_addr[5:0])
                6'd0  : o_data <= 64'h708898A8C8887000; // 0
                6'd1  : o_data <= 64'h2060202020207000; // 1
                6'd2  : o_data <= 64'h708808102040F800; // 2
                6'd3  : o_data <= 64'hF810201008887000; // 3
                6'd4  : o_data <= 64'h10305090F8101000; // 4
                6'd5  : o_data <= 64'hF880F00808887000; // 5
                6'd6  : o_data <= 64'h304080F088887000; // 6
                6'd7  : o_data <= 64'hF808102040404000; // 7
                6'd8  : o_data <= 64'h7088887088887000; // 8
                6'd9  : o_data <= 64'h7088887808106000; // 9
                6'd10 : o_data <= 64'h70888888F8888800; // A
                6'd11 : o_data <= 64'hF08888F08888F000; // B
                6'd12 : o_data <= 64'h7088808080887000; // C
                6'd13 : o_data <= 64'hE09088888890E000; // D
                6'd14 : o_data <= 64'hF88080F08080F800; // E
                6'd15 : o_data <= 64'hF88080F080808000; // F
                6'd16 : o_data <= 64'h708880B888887800; // G
                6'd17 : o_data <= 64'h888888F888888800; // H
                6'd18 : o_data <= 64'h7020202020207000; // I
                6'd19 : o_data <= 64'h3810101010906000; // J
                6'd20 : o_data <= 64'h8890A0C0A0908800; // K
                6'd21 : o_data <= 64'h808080808080F800; // L
                6'd22 : o_data <= 64'h88D8A8A888888800; // M
                6'd23 : o_data <= 64'h8888C8A898888800; // N
                6'd24 : o_data <= 64'h7088888888887000; // O
                6'd25 : o_data <= 64'hF08888F080808000; // P
                6'd26 : o_data <= 64'h70888888A8906800; // Q
                6'd27 : o_data <= 64'hF08888F0A0908800; // R
                6'd28 : o_data <= 64'h788080700808F000; // S
                6'd29 : o_data <= 64'hF820202020202000; // T
                6'd30 : o_data <= 64'h8888888888887000; // U
                6'd31 : o_data <= 64'h8888888888502000; // V
                6'd32 : o_data <= 64'h888888A8A8A85000; // W
                6'd33 : o_data <= 64'h8888502050888800; // X
                6'd34 : o_data <= 64'h8888502020202000; // Y
                6'd35 : o_data <= 64'hF80810204080F800; // Z
                6'd36 : o_data <= 64'h7040404040407000; // [
                6'd37 : o_data <= 64'h8850F820F8202000; // ¥
                6'd38 : o_data <= 64'h7010101010107000; // ]
                6'd39 : o_data <= 64'h2050880000000000; // ^
                6'd40 : o_data <= 64'h000000000000F800; // _
                6'd41 : o_data <= 64'h0060600060600000; // :
                6'd42 : o_data <= 64'h0000000000000000; // " "
                default : o_data <= 64'd0;
            endcase
        end
    end

endmodule

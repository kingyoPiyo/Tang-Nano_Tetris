/********************************************************
* Title    : BGM ROM (Korobushka)
* Date     : 2020/11/07
* Design   : kingyo
* Note     : o_data[31:15] : DeltaTime[ms]
             o_data[15: 8] : EventType
             o_data[ 7: 0] : Param1
********************************************************/
module bgm_rom (
    input   wire            i_clk,
    input   wire            i_res_n,
    input   wire    [ 9:0]  i_addr,
    output  reg     [31:0]  o_data
    )/* synthesis syn_romstyle = "block_rom" */;

    always @(posedge i_clk or negedge i_res_n) begin
        if (~i_res_n) begin
            o_data <= 32'd0;
        end else begin
            case (i_addr[9:0])
                10'd0: o_data <= 32'h00009128;
                10'd1: o_data <= 32'h00F09134;
                10'd2: o_data <= 32'h00F09128;
                10'd3: o_data <= 32'h00F09134;
                10'd4: o_data <= 32'h00F09128;
                10'd5: o_data <= 32'h00F09134;
                10'd6: o_data <= 32'h00F09128;
                10'd7: o_data <= 32'h00F09134;
                10'd8: o_data <= 32'h00F0912D;
                10'd9: o_data <= 32'h00F09139;
                10'd10: o_data <= 32'h00F0912D;
                10'd11: o_data <= 32'h00F09139;
                10'd12: o_data <= 32'h00F0912D;
                10'd13: o_data <= 32'h00F09139;
                10'd14: o_data <= 32'h00F0912D;
                10'd15: o_data <= 32'h00F09139;
                10'd16: o_data <= 32'h00F0904C;
                10'd17: o_data <= 32'h00009128;
                10'd18: o_data <= 32'h00F0804C;
                10'd19: o_data <= 32'h00009134;
                10'd20: o_data <= 32'h00F09047;
                10'd21: o_data <= 32'h00009128;
                10'd22: o_data <= 32'h00F08047;
                10'd23: o_data <= 32'h00009048;
                10'd24: o_data <= 32'h00009134;
                10'd25: o_data <= 32'h00F08048;
                10'd26: o_data <= 32'h0000904A;
                10'd27: o_data <= 32'h00009128;
                10'd28: o_data <= 32'h00F0804A;
                10'd29: o_data <= 32'h0000904C;
                10'd30: o_data <= 32'h00009134;
                10'd31: o_data <= 32'h0078804C;
                10'd32: o_data <= 32'h0000904A;
                10'd33: o_data <= 32'h0078804A;
                10'd34: o_data <= 32'h00009048;
                10'd35: o_data <= 32'h00009128;
                10'd36: o_data <= 32'h00F08048;
                10'd37: o_data <= 32'h00009047;
                10'd38: o_data <= 32'h00009134;
                10'd39: o_data <= 32'h00F08047;
                10'd40: o_data <= 32'h00009045;
                10'd41: o_data <= 32'h0000912D;
                10'd42: o_data <= 32'h00F08045;
                10'd43: o_data <= 32'h00009139;
                10'd44: o_data <= 32'h00F09045;
                10'd45: o_data <= 32'h0000912D;
                10'd46: o_data <= 32'h00F08045;
                10'd47: o_data <= 32'h00009048;
                10'd48: o_data <= 32'h00009139;
                10'd49: o_data <= 32'h00F08048;
                10'd50: o_data <= 32'h0000904C;
                10'd51: o_data <= 32'h0000912D;
                10'd52: o_data <= 32'h00F0804C;
                10'd53: o_data <= 32'h00009139;
                10'd54: o_data <= 32'h00F0904A;
                10'd55: o_data <= 32'h0000912D;
                10'd56: o_data <= 32'h00F0804A;
                10'd57: o_data <= 32'h00009048;
                10'd58: o_data <= 32'h00009139;
                10'd59: o_data <= 32'h00F08048;
                10'd60: o_data <= 32'h00009047;
                10'd61: o_data <= 32'h0000912C;
                10'd62: o_data <= 32'h00F08047;
                10'd63: o_data <= 32'h00009138;
                10'd64: o_data <= 32'h00F08138;
                10'd65: o_data <= 32'h0000912C;
                10'd66: o_data <= 32'h00F09048;
                10'd67: o_data <= 32'h00009138;
                10'd68: o_data <= 32'h00F08048;
                10'd69: o_data <= 32'h0000904A;
                10'd70: o_data <= 32'h00009128;
                10'd71: o_data <= 32'h00F0804A;
                10'd72: o_data <= 32'h00009134;
                10'd73: o_data <= 32'h00F0904C;
                10'd74: o_data <= 32'h00009128;
                10'd75: o_data <= 32'h00F0804C;
                10'd76: o_data <= 32'h00009134;
                10'd77: o_data <= 32'h00F09048;
                10'd78: o_data <= 32'h0000912D;
                10'd79: o_data <= 32'h00F08048;
                10'd80: o_data <= 32'h00009139;
                10'd81: o_data <= 32'h00F09045;
                10'd82: o_data <= 32'h0000912D;
                10'd83: o_data <= 32'h00F08045;
                10'd84: o_data <= 32'h00009139;
                10'd85: o_data <= 32'h00F09045;
                10'd86: o_data <= 32'h0000912D;
                10'd87: o_data <= 32'h00F08045;
                10'd88: o_data <= 32'h00009139;
                10'd89: o_data <= 32'h00F08139;
                10'd90: o_data <= 32'h0000912F;
                10'd91: o_data <= 32'h00F0812F;
                10'd92: o_data <= 32'h00009130;
                10'd93: o_data <= 32'h00F08130;
                10'd94: o_data <= 32'h00009132;
                10'd95: o_data <= 32'h00F0904A;
                10'd96: o_data <= 32'h00009126;
                10'd97: o_data <= 32'h00F0804A;
                10'd98: o_data <= 32'h00008126;
                10'd99: o_data <= 32'h00F0904D;
                10'd100: o_data <= 32'h00009126;
                10'd101: o_data <= 32'h00F0804D;
                10'd102: o_data <= 32'h00009051;
                10'd103: o_data <= 32'h00008126;
                10'd104: o_data <= 32'h00F08051;
                10'd105: o_data <= 32'h00009126;
                10'd106: o_data <= 32'h00788126;
                10'd107: o_data <= 32'h00009126;
                10'd108: o_data <= 32'h0078904F;
                10'd109: o_data <= 32'h0000912D;
                10'd110: o_data <= 32'h00F0804F;
                10'd111: o_data <= 32'h0000904D;
                10'd112: o_data <= 32'h0000912B;
                10'd113: o_data <= 32'h00F0804D;
                10'd114: o_data <= 32'h0000904C;
                10'd115: o_data <= 32'h00009124;
                10'd116: o_data <= 32'h00F0804C;
                10'd117: o_data <= 32'h00009130;
                10'd118: o_data <= 32'h00F08130;
                10'd119: o_data <= 32'h00009124;
                10'd120: o_data <= 32'h00F09048;
                10'd121: o_data <= 32'h00009130;
                10'd122: o_data <= 32'h00F08048;
                10'd123: o_data <= 32'h0000904C;
                10'd124: o_data <= 32'h00009124;
                10'd125: o_data <= 32'h00F0804C;
                10'd126: o_data <= 32'h0000904D;
                10'd127: o_data <= 32'h0000912B;
                10'd128: o_data <= 32'h0078804D;
                10'd129: o_data <= 32'h0000904C;
                10'd130: o_data <= 32'h0078804C;
                10'd131: o_data <= 32'h0000904A;
                10'd132: o_data <= 32'h00009124;
                10'd133: o_data <= 32'h00F0804A;
                10'd134: o_data <= 32'h00009048;
                10'd135: o_data <= 32'h0000912B;
                10'd136: o_data <= 32'h00F08048;
                10'd137: o_data <= 32'h00009047;
                10'd138: o_data <= 32'h0000912F;
                10'd139: o_data <= 32'h00F08047;
                10'd140: o_data <= 32'h0000913B;
                10'd141: o_data <= 32'h00F0813B;
                10'd142: o_data <= 32'h00F09048;
                10'd143: o_data <= 32'h0000913B;
                10'd144: o_data <= 32'h00F08048;
                10'd145: o_data <= 32'h0000904A;
                10'd146: o_data <= 32'h00009134;
                10'd147: o_data <= 32'h00F0804A;
                10'd148: o_data <= 32'h00009044;
                10'd149: o_data <= 32'h00008134;
                10'd150: o_data <= 32'h00F08044;
                10'd151: o_data <= 32'h0000904C;
                10'd152: o_data <= 32'h00009138;
                10'd153: o_data <= 32'h00F0804C;
                10'd154: o_data <= 32'h00009044;
                10'd155: o_data <= 32'h00008138;
                10'd156: o_data <= 32'h00F08044;
                10'd157: o_data <= 32'h00009048;
                10'd158: o_data <= 32'h0000912D;
                10'd159: o_data <= 32'h00F08048;
                10'd160: o_data <= 32'h00009134;
                10'd161: o_data <= 32'h00F09045;
                10'd162: o_data <= 32'h0000912D;
                10'd163: o_data <= 32'h00F08045;
                10'd164: o_data <= 32'h00009134;
                10'd165: o_data <= 32'h00F09045;
                10'd166: o_data <= 32'h0000912D;
                10'd167: o_data <= 32'h00F0812D;
                10'd168: o_data <= 32'h00009134;
                10'd169: o_data <= 32'h00F08134;
                10'd170: o_data <= 32'h00009134;
                10'd171: o_data <= 32'h00F08134;
                10'd172: o_data <= 32'h00009134;
                10'd173: o_data <= 32'h00F08045;
                10'd174: o_data <= 32'h0000904C;
                10'd175: o_data <= 32'h00009128;
                10'd176: o_data <= 32'h00F0804C;
                10'd177: o_data <= 32'h00009134;
                10'd178: o_data <= 32'h00F09047;
                10'd179: o_data <= 32'h00009128;
                10'd180: o_data <= 32'h00F08047;
                10'd181: o_data <= 32'h00009048;
                10'd182: o_data <= 32'h00009134;
                10'd183: o_data <= 32'h00F08048;
                10'd184: o_data <= 32'h0000904A;
                10'd185: o_data <= 32'h00009128;
                10'd186: o_data <= 32'h00F0804A;
                10'd187: o_data <= 32'h0000904C;
                10'd188: o_data <= 32'h00009134;
                10'd189: o_data <= 32'h0078804C;
                10'd190: o_data <= 32'h0000904A;
                10'd191: o_data <= 32'h0078804A;
                10'd192: o_data <= 32'h00009048;
                10'd193: o_data <= 32'h00009128;
                10'd194: o_data <= 32'h00F08048;
                10'd195: o_data <= 32'h00009047;
                10'd196: o_data <= 32'h00009134;
                10'd197: o_data <= 32'h00F08047;
                10'd198: o_data <= 32'h00009045;
                10'd199: o_data <= 32'h0000912D;
                10'd200: o_data <= 32'h00F08045;
                10'd201: o_data <= 32'h00009139;
                10'd202: o_data <= 32'h00F09045;
                10'd203: o_data <= 32'h0000912D;
                10'd204: o_data <= 32'h00F08045;
                10'd205: o_data <= 32'h00009048;
                10'd206: o_data <= 32'h00009139;
                10'd207: o_data <= 32'h00F08048;
                10'd208: o_data <= 32'h0000904C;
                10'd209: o_data <= 32'h0000912D;
                10'd210: o_data <= 32'h00F0804C;
                10'd211: o_data <= 32'h00009139;
                10'd212: o_data <= 32'h00F0904A;
                10'd213: o_data <= 32'h0000912D;
                10'd214: o_data <= 32'h00F0804A;
                10'd215: o_data <= 32'h00009048;
                10'd216: o_data <= 32'h00009139;
                10'd217: o_data <= 32'h00F08048;
                10'd218: o_data <= 32'h00009047;
                10'd219: o_data <= 32'h0000912C;
                10'd220: o_data <= 32'h00F08047;
                10'd221: o_data <= 32'h00009138;
                10'd222: o_data <= 32'h00F08138;
                10'd223: o_data <= 32'h0000912C;
                10'd224: o_data <= 32'h00F09048;
                10'd225: o_data <= 32'h00009138;
                10'd226: o_data <= 32'h00F08048;
                10'd227: o_data <= 32'h0000904A;
                10'd228: o_data <= 32'h00009128;
                10'd229: o_data <= 32'h00F0804A;
                10'd230: o_data <= 32'h00009134;
                10'd231: o_data <= 32'h00F0904C;
                10'd232: o_data <= 32'h00009128;
                10'd233: o_data <= 32'h00F0804C;
                10'd234: o_data <= 32'h00009134;
                10'd235: o_data <= 32'h00F09048;
                10'd236: o_data <= 32'h0000912D;
                10'd237: o_data <= 32'h00F08048;
                10'd238: o_data <= 32'h00009139;
                10'd239: o_data <= 32'h00F09045;
                10'd240: o_data <= 32'h0000912D;
                10'd241: o_data <= 32'h00F08045;
                10'd242: o_data <= 32'h00009139;
                10'd243: o_data <= 32'h00F09045;
                10'd244: o_data <= 32'h0000912D;
                10'd245: o_data <= 32'h00F08045;
                10'd246: o_data <= 32'h00009139;
                10'd247: o_data <= 32'h00F08139;
                10'd248: o_data <= 32'h0000912F;
                10'd249: o_data <= 32'h00F0812F;
                10'd250: o_data <= 32'h00009130;
                10'd251: o_data <= 32'h00F08130;
                10'd252: o_data <= 32'h00009132;
                10'd253: o_data <= 32'h00F0904A;
                10'd254: o_data <= 32'h00009126;
                10'd255: o_data <= 32'h00F0804A;
                10'd256: o_data <= 32'h00008126;
                10'd257: o_data <= 32'h00F0904D;
                10'd258: o_data <= 32'h00009126;
                10'd259: o_data <= 32'h00F0804D;
                10'd260: o_data <= 32'h00009051;
                10'd261: o_data <= 32'h00008126;
                10'd262: o_data <= 32'h00F08051;
                10'd263: o_data <= 32'h00009126;
                10'd264: o_data <= 32'h00788126;
                10'd265: o_data <= 32'h00009126;
                10'd266: o_data <= 32'h0078904F;
                10'd267: o_data <= 32'h0000912D;
                10'd268: o_data <= 32'h00F0804F;
                10'd269: o_data <= 32'h0000904D;
                10'd270: o_data <= 32'h0000912B;
                10'd271: o_data <= 32'h00F0804D;
                10'd272: o_data <= 32'h0000904C;
                10'd273: o_data <= 32'h00009124;
                10'd274: o_data <= 32'h00F0804C;
                10'd275: o_data <= 32'h00009130;
                10'd276: o_data <= 32'h00F08130;
                10'd277: o_data <= 32'h00009124;
                10'd278: o_data <= 32'h00F09048;
                10'd279: o_data <= 32'h00009130;
                10'd280: o_data <= 32'h00F08048;
                10'd281: o_data <= 32'h0000904C;
                10'd282: o_data <= 32'h00009124;
                10'd283: o_data <= 32'h00F0804C;
                10'd284: o_data <= 32'h0000904D;
                10'd285: o_data <= 32'h0000912B;
                10'd286: o_data <= 32'h0078804D;
                10'd287: o_data <= 32'h0000904C;
                10'd288: o_data <= 32'h0078804C;
                10'd289: o_data <= 32'h0000904A;
                10'd290: o_data <= 32'h00009124;
                10'd291: o_data <= 32'h00F0804A;
                10'd292: o_data <= 32'h00009048;
                10'd293: o_data <= 32'h0000912B;
                10'd294: o_data <= 32'h00F08048;
                10'd295: o_data <= 32'h00009047;
                10'd296: o_data <= 32'h0000912F;
                10'd297: o_data <= 32'h00F08047;
                10'd298: o_data <= 32'h0000913B;
                10'd299: o_data <= 32'h00F0813B;
                10'd300: o_data <= 32'h00F09048;
                10'd301: o_data <= 32'h0000913B;
                10'd302: o_data <= 32'h00F08048;
                10'd303: o_data <= 32'h0000904A;
                10'd304: o_data <= 32'h00009134;
                10'd305: o_data <= 32'h00F0804A;
                10'd306: o_data <= 32'h00009044;
                10'd307: o_data <= 32'h00008134;
                10'd308: o_data <= 32'h00F08044;
                10'd309: o_data <= 32'h0000904C;
                10'd310: o_data <= 32'h00009138;
                10'd311: o_data <= 32'h00F0804C;
                10'd312: o_data <= 32'h00009044;
                10'd313: o_data <= 32'h00008138;
                10'd314: o_data <= 32'h00F08044;
                10'd315: o_data <= 32'h00009048;
                10'd316: o_data <= 32'h0000912D;
                10'd317: o_data <= 32'h00F08048;
                10'd318: o_data <= 32'h00009134;
                10'd319: o_data <= 32'h00F09045;
                10'd320: o_data <= 32'h0000912D;
                10'd321: o_data <= 32'h00F08045;
                10'd322: o_data <= 32'h00009134;
                10'd323: o_data <= 32'h00F09045;
                10'd324: o_data <= 32'h0000912D;
                10'd325: o_data <= 32'h00F0812D;
                10'd326: o_data <= 32'h00009134;
                10'd327: o_data <= 32'h00F08134;
                10'd328: o_data <= 32'h00009134;
                10'd329: o_data <= 32'h00F08134;
                10'd330: o_data <= 32'h00009134;
                10'd331: o_data <= 32'h00F08045;
                10'd332: o_data <= 32'h00009040;
                10'd333: o_data <= 32'h0000912D;
                10'd334: o_data <= 32'h00F0812D;
                10'd335: o_data <= 32'h00009134;
                10'd336: o_data <= 32'h00F08134;
                10'd337: o_data <= 32'h0000912D;
                10'd338: o_data <= 32'h00F0812D;
                10'd339: o_data <= 32'h00009134;
                10'd340: o_data <= 32'h00F08040;
                10'd341: o_data <= 32'h0000903C;
                10'd342: o_data <= 32'h0000912D;
                10'd343: o_data <= 32'h00F0812D;
                10'd344: o_data <= 32'h00009134;
                10'd345: o_data <= 32'h00F08134;
                10'd346: o_data <= 32'h0000912D;
                10'd347: o_data <= 32'h00F0812D;
                10'd348: o_data <= 32'h00009134;
                10'd349: o_data <= 32'h00F0803C;
                10'd350: o_data <= 32'h0000903E;
                10'd351: o_data <= 32'h0000912C;
                10'd352: o_data <= 32'h00F0812C;
                10'd353: o_data <= 32'h00009134;
                10'd354: o_data <= 32'h00F08134;
                10'd355: o_data <= 32'h0000912C;
                10'd356: o_data <= 32'h00F0812C;
                10'd357: o_data <= 32'h00009134;
                10'd358: o_data <= 32'h00F0803E;
                10'd359: o_data <= 32'h0000903B;
                10'd360: o_data <= 32'h0000912C;
                10'd361: o_data <= 32'h00F0812C;
                10'd362: o_data <= 32'h00009134;
                10'd363: o_data <= 32'h00F08134;
                10'd364: o_data <= 32'h0000912C;
                10'd365: o_data <= 32'h00F0812C;
                10'd366: o_data <= 32'h00009134;
                10'd367: o_data <= 32'h00F0803B;
                10'd368: o_data <= 32'h0000903C;
                10'd369: o_data <= 32'h0000912D;
                10'd370: o_data <= 32'h00F0812D;
                10'd371: o_data <= 32'h00009134;
                10'd372: o_data <= 32'h00F08134;
                10'd373: o_data <= 32'h0000912D;
                10'd374: o_data <= 32'h00F0812D;
                10'd375: o_data <= 32'h00009134;
                10'd376: o_data <= 32'h00F0803C;
                10'd377: o_data <= 32'h00009039;
                10'd378: o_data <= 32'h0000912D;
                10'd379: o_data <= 32'h00F0812D;
                10'd380: o_data <= 32'h00009134;
                10'd381: o_data <= 32'h00F08134;
                10'd382: o_data <= 32'h0000912D;
                10'd383: o_data <= 32'h00F0812D;
                10'd384: o_data <= 32'h00009134;
                10'd385: o_data <= 32'h00F08039;
                10'd386: o_data <= 32'h00009038;
                10'd387: o_data <= 32'h0000912C;
                10'd388: o_data <= 32'h00F0812C;
                10'd389: o_data <= 32'h00009134;
                10'd390: o_data <= 32'h00F08134;
                10'd391: o_data <= 32'h0000912C;
                10'd392: o_data <= 32'h00F0812C;
                10'd393: o_data <= 32'h00009134;
                10'd394: o_data <= 32'h00F08038;
                10'd395: o_data <= 32'h0000903B;
                10'd396: o_data <= 32'h0000912C;
                10'd397: o_data <= 32'h00F0812C;
                10'd398: o_data <= 32'h00009134;
                10'd399: o_data <= 32'h00F08134;
                10'd400: o_data <= 32'h0000912C;
                10'd401: o_data <= 32'h00F0812C;
                10'd402: o_data <= 32'h00009134;
                10'd403: o_data <= 32'h00F0803B;
                10'd404: o_data <= 32'h00009040;
                10'd405: o_data <= 32'h0000912D;
                10'd406: o_data <= 32'h00F0812D;
                10'd407: o_data <= 32'h00009134;
                10'd408: o_data <= 32'h00F08134;
                10'd409: o_data <= 32'h0000912D;
                10'd410: o_data <= 32'h00F0812D;
                10'd411: o_data <= 32'h00009134;
                10'd412: o_data <= 32'h00F08040;
                10'd413: o_data <= 32'h0000903C;
                10'd414: o_data <= 32'h0000912D;
                10'd415: o_data <= 32'h00F0812D;
                10'd416: o_data <= 32'h00009134;
                10'd417: o_data <= 32'h00F08134;
                10'd418: o_data <= 32'h0000912D;
                10'd419: o_data <= 32'h00F0812D;
                10'd420: o_data <= 32'h00009134;
                10'd421: o_data <= 32'h00F0803C;
                10'd422: o_data <= 32'h0000903E;
                10'd423: o_data <= 32'h0000912C;
                10'd424: o_data <= 32'h00F0812C;
                10'd425: o_data <= 32'h00009134;
                10'd426: o_data <= 32'h00F08134;
                10'd427: o_data <= 32'h0000912C;
                10'd428: o_data <= 32'h00F0812C;
                10'd429: o_data <= 32'h00009134;
                10'd430: o_data <= 32'h00F0803E;
                10'd431: o_data <= 32'h0000903B;
                10'd432: o_data <= 32'h0000912C;
                10'd433: o_data <= 32'h00F0812C;
                10'd434: o_data <= 32'h00009134;
                10'd435: o_data <= 32'h00F08134;
                10'd436: o_data <= 32'h0000912C;
                10'd437: o_data <= 32'h00F0812C;
                10'd438: o_data <= 32'h00009134;
                10'd439: o_data <= 32'h00F0803B;
                10'd440: o_data <= 32'h0000903C;
                10'd441: o_data <= 32'h0000912D;
                10'd442: o_data <= 32'h00F0812D;
                10'd443: o_data <= 32'h00009134;
                10'd444: o_data <= 32'h00F0803C;
                10'd445: o_data <= 32'h00009040;
                10'd446: o_data <= 32'h0000912D;
                10'd447: o_data <= 32'h00F0812D;
                10'd448: o_data <= 32'h00009134;
                10'd449: o_data <= 32'h00F08040;
                10'd450: o_data <= 32'h00009045;
                10'd451: o_data <= 32'h0000912D;
                10'd452: o_data <= 32'h00F0812D;
                10'd453: o_data <= 32'h00009134;
                10'd454: o_data <= 32'h00F08134;
                10'd455: o_data <= 32'h0000912D;
                10'd456: o_data <= 32'h00F0812D;
                10'd457: o_data <= 32'h00009134;
                10'd458: o_data <= 32'h00F08045;
                10'd459: o_data <= 32'h00009044;
                10'd460: o_data <= 32'h0000912C;
                10'd461: o_data <= 32'h00F0812C;
                10'd462: o_data <= 32'h00009134;
                10'd463: o_data <= 32'h00F08134;
                10'd464: o_data <= 32'h0000912C;
                10'd465: o_data <= 32'h00F0812C;
                10'd466: o_data <= 32'h00009134;
                10'd467: o_data <= 32'h00F08134;
                10'd468: o_data <= 32'h0000912C;
                10'd469: o_data <= 32'h00F0812C;
                10'd470: o_data <= 32'h00009134;
                10'd471: o_data <= 32'h00F08134;
                10'd472: o_data <= 32'h0000912C;
                10'd473: o_data <= 32'h00F0812C;
                10'd474: o_data <= 32'h00009134;
                10'd475: o_data <= 32'h00F08044;
                10'd476: o_data <= 32'h0000904C;
                10'd477: o_data <= 32'h00009128;
                10'd478: o_data <= 32'h00F0804C;
                10'd479: o_data <= 32'h00009134;
                10'd480: o_data <= 32'h00F09047;
                10'd481: o_data <= 32'h00009128;
                10'd482: o_data <= 32'h00F08047;
                10'd483: o_data <= 32'h00009048;
                10'd484: o_data <= 32'h00009134;
                10'd485: o_data <= 32'h00F08048;
                10'd486: o_data <= 32'h0000904A;
                10'd487: o_data <= 32'h00009128;
                10'd488: o_data <= 32'h00F0804A;
                10'd489: o_data <= 32'h0000904C;
                10'd490: o_data <= 32'h00009134;
                10'd491: o_data <= 32'h0078804C;
                10'd492: o_data <= 32'h0000904A;
                10'd493: o_data <= 32'h0078804A;
                10'd494: o_data <= 32'h00009048;
                10'd495: o_data <= 32'h00009128;
                10'd496: o_data <= 32'h00F08048;
                10'd497: o_data <= 32'h00009047;
                10'd498: o_data <= 32'h00009134;
                10'd499: o_data <= 32'h00F08047;
                10'd500: o_data <= 32'h00009045;
                10'd501: o_data <= 32'h0000912D;
                10'd502: o_data <= 32'h00F08045;
                10'd503: o_data <= 32'h00009139;
                10'd504: o_data <= 32'h00F09045;
                10'd505: o_data <= 32'h0000912D;
                10'd506: o_data <= 32'h00F08045;
                10'd507: o_data <= 32'h00009048;
                10'd508: o_data <= 32'h00009139;
                10'd509: o_data <= 32'h00F08048;
                10'd510: o_data <= 32'h0000904C;
                10'd511: o_data <= 32'h0000912D;
                10'd512: o_data <= 32'h00F0804C;
                10'd513: o_data <= 32'h00009139;
                10'd514: o_data <= 32'h00F0904A;
                10'd515: o_data <= 32'h0000912D;
                10'd516: o_data <= 32'h00F0804A;
                10'd517: o_data <= 32'h00009048;
                10'd518: o_data <= 32'h00009139;
                10'd519: o_data <= 32'h00F08048;
                10'd520: o_data <= 32'h00009047;
                10'd521: o_data <= 32'h0000912C;
                10'd522: o_data <= 32'h00F08047;
                10'd523: o_data <= 32'h00009138;
                10'd524: o_data <= 32'h00F08138;
                10'd525: o_data <= 32'h0000912C;
                10'd526: o_data <= 32'h00F09048;
                10'd527: o_data <= 32'h00009138;
                10'd528: o_data <= 32'h00F08048;
                10'd529: o_data <= 32'h0000904A;
                10'd530: o_data <= 32'h00009128;
                10'd531: o_data <= 32'h00F0804A;
                10'd532: o_data <= 32'h00009134;
                10'd533: o_data <= 32'h00F0904C;
                10'd534: o_data <= 32'h00009128;
                10'd535: o_data <= 32'h00F0804C;
                10'd536: o_data <= 32'h00009134;
                10'd537: o_data <= 32'h00F09048;
                10'd538: o_data <= 32'h0000912D;
                10'd539: o_data <= 32'h00F08048;
                10'd540: o_data <= 32'h00009139;
                10'd541: o_data <= 32'h00F09045;
                10'd542: o_data <= 32'h0000912D;
                10'd543: o_data <= 32'h00F08045;
                10'd544: o_data <= 32'h00009139;
                10'd545: o_data <= 32'h00F09045;
                10'd546: o_data <= 32'h0000912D;
                10'd547: o_data <= 32'h00F08045;
                10'd548: o_data <= 32'h00009139;
                10'd549: o_data <= 32'h00F08139;
                10'd550: o_data <= 32'h0000912F;
                10'd551: o_data <= 32'h00F0812F;
                10'd552: o_data <= 32'h00009130;
                10'd553: o_data <= 32'h00F08130;
                10'd554: o_data <= 32'h00009132;
                10'd555: o_data <= 32'h00F0904A;
                10'd556: o_data <= 32'h00009126;
                10'd557: o_data <= 32'h00F0804A;
                10'd558: o_data <= 32'h00008126;
                10'd559: o_data <= 32'h00F0904D;
                10'd560: o_data <= 32'h00009126;
                10'd561: o_data <= 32'h00F0804D;
                10'd562: o_data <= 32'h00009051;
                10'd563: o_data <= 32'h00008126;
                10'd564: o_data <= 32'h00F08051;
                10'd565: o_data <= 32'h00009126;
                10'd566: o_data <= 32'h00788126;
                10'd567: o_data <= 32'h00009126;
                10'd568: o_data <= 32'h0078904F;
                10'd569: o_data <= 32'h0000912D;
                10'd570: o_data <= 32'h00F0804F;
                10'd571: o_data <= 32'h0000904D;
                10'd572: o_data <= 32'h0000912B;
                10'd573: o_data <= 32'h00F0804D;
                10'd574: o_data <= 32'h0000904C;
                10'd575: o_data <= 32'h00009124;
                10'd576: o_data <= 32'h00F0804C;
                10'd577: o_data <= 32'h00009130;
                10'd578: o_data <= 32'h00F08130;
                10'd579: o_data <= 32'h00009124;
                10'd580: o_data <= 32'h00F09048;
                10'd581: o_data <= 32'h00009130;
                10'd582: o_data <= 32'h00F08048;
                10'd583: o_data <= 32'h0000904C;
                10'd584: o_data <= 32'h00009124;
                10'd585: o_data <= 32'h00F0804C;
                10'd586: o_data <= 32'h0000904D;
                10'd587: o_data <= 32'h0000912B;
                10'd588: o_data <= 32'h0078804D;
                10'd589: o_data <= 32'h0000904C;
                10'd590: o_data <= 32'h0078804C;
                10'd591: o_data <= 32'h0000904A;
                10'd592: o_data <= 32'h00009124;
                10'd593: o_data <= 32'h00F0804A;
                10'd594: o_data <= 32'h00009048;
                10'd595: o_data <= 32'h0000912B;
                10'd596: o_data <= 32'h00F08048;
                10'd597: o_data <= 32'h00009047;
                10'd598: o_data <= 32'h0000912F;
                10'd599: o_data <= 32'h00F08047;
                10'd600: o_data <= 32'h0000913B;
                10'd601: o_data <= 32'h00F0813B;
                10'd602: o_data <= 32'h00F09048;
                10'd603: o_data <= 32'h0000913B;
                10'd604: o_data <= 32'h00F08048;
                10'd605: o_data <= 32'h0000904A;
                10'd606: o_data <= 32'h00009134;
                10'd607: o_data <= 32'h00F0804A;
                10'd608: o_data <= 32'h00009044;
                10'd609: o_data <= 32'h00008134;
                10'd610: o_data <= 32'h00F08044;
                10'd611: o_data <= 32'h0000904C;
                10'd612: o_data <= 32'h00009138;
                10'd613: o_data <= 32'h00F0804C;
                10'd614: o_data <= 32'h00009044;
                10'd615: o_data <= 32'h00008138;
                10'd616: o_data <= 32'h00F08044;
                10'd617: o_data <= 32'h00009048;
                10'd618: o_data <= 32'h0000912D;
                10'd619: o_data <= 32'h00F08048;
                10'd620: o_data <= 32'h00009134;
                10'd621: o_data <= 32'h00F09045;
                10'd622: o_data <= 32'h0000912D;
                10'd623: o_data <= 32'h00F08045;
                10'd624: o_data <= 32'h00009134;
                10'd625: o_data <= 32'h00F09045;
                10'd626: o_data <= 32'h0000912D;
                10'd627: o_data <= 32'h03C08045;
                10'd628: o_data <= 32'h0000904C;
                10'd629: o_data <= 32'h00009128;
                10'd630: o_data <= 32'h00F0804C;
                10'd631: o_data <= 32'h00009134;
                10'd632: o_data <= 32'h00F09047;
                10'd633: o_data <= 32'h00009128;
                10'd634: o_data <= 32'h00F08047;
                10'd635: o_data <= 32'h00009048;
                10'd636: o_data <= 32'h00009134;
                10'd637: o_data <= 32'h00F08048;
                10'd638: o_data <= 32'h0000904A;
                10'd639: o_data <= 32'h00009128;
                10'd640: o_data <= 32'h00F0804A;
                10'd641: o_data <= 32'h0000904C;
                10'd642: o_data <= 32'h00009134;
                10'd643: o_data <= 32'h0078804C;
                10'd644: o_data <= 32'h0000904A;
                10'd645: o_data <= 32'h0078804A;
                10'd646: o_data <= 32'h00009048;
                10'd647: o_data <= 32'h00009128;
                10'd648: o_data <= 32'h00F08048;
                10'd649: o_data <= 32'h00009047;
                10'd650: o_data <= 32'h00009134;
                10'd651: o_data <= 32'h00F08047;
                10'd652: o_data <= 32'h00009045;
                10'd653: o_data <= 32'h0000912D;
                10'd654: o_data <= 32'h00F08045;
                10'd655: o_data <= 32'h00009139;
                10'd656: o_data <= 32'h00F09045;
                10'd657: o_data <= 32'h0000912D;
                10'd658: o_data <= 32'h00F08045;
                10'd659: o_data <= 32'h00009048;
                10'd660: o_data <= 32'h00009139;
                10'd661: o_data <= 32'h00F08048;
                10'd662: o_data <= 32'h0000904C;
                10'd663: o_data <= 32'h0000912D;
                10'd664: o_data <= 32'h00F0804C;
                10'd665: o_data <= 32'h00009139;
                10'd666: o_data <= 32'h00F0904A;
                10'd667: o_data <= 32'h0000912D;
                10'd668: o_data <= 32'h00F0804A;
                10'd669: o_data <= 32'h00009048;
                10'd670: o_data <= 32'h00009139;
                10'd671: o_data <= 32'h00F08048;
                10'd672: o_data <= 32'h00009047;
                10'd673: o_data <= 32'h0000912C;
                10'd674: o_data <= 32'h00F08047;
                10'd675: o_data <= 32'h00009138;
                10'd676: o_data <= 32'h00F08138;
                10'd677: o_data <= 32'h0000912C;
                10'd678: o_data <= 32'h00F09048;
                10'd679: o_data <= 32'h00009138;
                10'd680: o_data <= 32'h00F08048;
                10'd681: o_data <= 32'h0000904A;
                10'd682: o_data <= 32'h00009128;
                10'd683: o_data <= 32'h00F0804A;
                10'd684: o_data <= 32'h00009134;
                10'd685: o_data <= 32'h00F0904C;
                10'd686: o_data <= 32'h00009128;
                10'd687: o_data <= 32'h00F0804C;
                10'd688: o_data <= 32'h00009134;
                10'd689: o_data <= 32'h00F09048;
                10'd690: o_data <= 32'h0000912D;
                10'd691: o_data <= 32'h00F08048;
                10'd692: o_data <= 32'h00009139;
                10'd693: o_data <= 32'h00F09045;
                10'd694: o_data <= 32'h0000912D;
                10'd695: o_data <= 32'h00F08045;
                10'd696: o_data <= 32'h00009139;
                10'd697: o_data <= 32'h00F09045;
                10'd698: o_data <= 32'h0000912D;
                10'd699: o_data <= 32'h00F08045;
                10'd700: o_data <= 32'h00009139;
                10'd701: o_data <= 32'h00F08139;
                10'd702: o_data <= 32'h0000912F;
                10'd703: o_data <= 32'h00F0812F;
                10'd704: o_data <= 32'h00009130;
                10'd705: o_data <= 32'h00F08130;
                10'd706: o_data <= 32'h00009132;
                10'd707: o_data <= 32'h00F0904A;
                10'd708: o_data <= 32'h00009126;
                10'd709: o_data <= 32'h00F0804A;
                10'd710: o_data <= 32'h00008126;
                10'd711: o_data <= 32'h00F0904D;
                10'd712: o_data <= 32'h00009126;
                10'd713: o_data <= 32'h00F0804D;
                10'd714: o_data <= 32'h00009051;
                10'd715: o_data <= 32'h00008126;
                10'd716: o_data <= 32'h00F08051;
                10'd717: o_data <= 32'h00009126;
                10'd718: o_data <= 32'h00788126;
                10'd719: o_data <= 32'h00009126;
                10'd720: o_data <= 32'h0078904F;
                10'd721: o_data <= 32'h0000912D;
                10'd722: o_data <= 32'h00F0804F;
                10'd723: o_data <= 32'h0000904D;
                10'd724: o_data <= 32'h0000912B;
                10'd725: o_data <= 32'h00F0804D;
                10'd726: o_data <= 32'h0000904C;
                10'd727: o_data <= 32'h00009124;
                10'd728: o_data <= 32'h00F0804C;
                10'd729: o_data <= 32'h00009130;
                10'd730: o_data <= 32'h00F08130;
                10'd731: o_data <= 32'h00009124;
                10'd732: o_data <= 32'h00F09048;
                10'd733: o_data <= 32'h00009130;
                10'd734: o_data <= 32'h00F08048;
                10'd735: o_data <= 32'h0000904C;
                10'd736: o_data <= 32'h00009124;
                10'd737: o_data <= 32'h00F0804C;
                10'd738: o_data <= 32'h0000904D;
                10'd739: o_data <= 32'h0000912B;
                10'd740: o_data <= 32'h0078804D;
                10'd741: o_data <= 32'h0000904C;
                10'd742: o_data <= 32'h0078804C;
                10'd743: o_data <= 32'h0000904A;
                10'd744: o_data <= 32'h00009124;
                10'd745: o_data <= 32'h00F0804A;
                10'd746: o_data <= 32'h00009048;
                10'd747: o_data <= 32'h0000912B;
                10'd748: o_data <= 32'h00F08048;
                10'd749: o_data <= 32'h00009047;
                10'd750: o_data <= 32'h0000912F;
                10'd751: o_data <= 32'h00F08047;
                10'd752: o_data <= 32'h0000913B;
                10'd753: o_data <= 32'h00F0813B;
                10'd754: o_data <= 32'h00F09048;
                10'd755: o_data <= 32'h0000913B;
                10'd756: o_data <= 32'h00F08048;
                10'd757: o_data <= 32'h0000904A;
                10'd758: o_data <= 32'h00009134;
                10'd759: o_data <= 32'h00F0804A;
                10'd760: o_data <= 32'h00009044;
                10'd761: o_data <= 32'h00008134;
                10'd762: o_data <= 32'h00F08044;
                10'd763: o_data <= 32'h0000904C;
                10'd764: o_data <= 32'h00009138;
                10'd765: o_data <= 32'h00F0804C;
                10'd766: o_data <= 32'h00009044;
                10'd767: o_data <= 32'h00008138;
                10'd768: o_data <= 32'h00F08044;
                10'd769: o_data <= 32'h00009048;
                10'd770: o_data <= 32'h0000912D;
                10'd771: o_data <= 32'h00F08048;
                10'd772: o_data <= 32'h00009134;
                10'd773: o_data <= 32'h00F09045;
                10'd774: o_data <= 32'h0000912D;
                10'd775: o_data <= 32'h00F08045;
                10'd776: o_data <= 32'h00009134;
                10'd777: o_data <= 32'h00F09045;
                10'd778: o_data <= 32'h0000912D;
                10'd779: o_data <= 32'h00F0812D;
                10'd780: o_data <= 32'h00009134;
                10'd781: o_data <= 32'h00F08134;
                10'd782: o_data <= 32'h00009134;
                10'd783: o_data <= 32'h00F08134;
                10'd784: o_data <= 32'h00009134;
                10'd785: o_data <= 32'h00F08045;
                10'd786: o_data <= 32'h0000904D;
                10'd787: o_data <= 32'h00009129;
                10'd788: o_data <= 32'h00F0804D;
                10'd789: o_data <= 32'h00009135;
                10'd790: o_data <= 32'h00F09048;
                10'd791: o_data <= 32'h00009129;
                10'd792: o_data <= 32'h00F08048;
                10'd793: o_data <= 32'h00009049;
                10'd794: o_data <= 32'h00009135;
                10'd795: o_data <= 32'h00F08049;
                10'd796: o_data <= 32'h0000904B;
                10'd797: o_data <= 32'h00009129;
                10'd798: o_data <= 32'h00F0804B;
                10'd799: o_data <= 32'h0000904D;
                10'd800: o_data <= 32'h00009135;
                10'd801: o_data <= 32'h0078804D;
                10'd802: o_data <= 32'h0000904B;
                10'd803: o_data <= 32'h0078804B;
                10'd804: o_data <= 32'h00009049;
                10'd805: o_data <= 32'h00009129;
                10'd806: o_data <= 32'h00F08049;
                10'd807: o_data <= 32'h00009048;
                10'd808: o_data <= 32'h00009135;
                10'd809: o_data <= 32'h00F08048;
                10'd810: o_data <= 32'h00009046;
                10'd811: o_data <= 32'h0000912E;
                10'd812: o_data <= 32'h00F08046;
                10'd813: o_data <= 32'h0000913A;
                10'd814: o_data <= 32'h00F09046;
                10'd815: o_data <= 32'h0000912E;
                10'd816: o_data <= 32'h00F08046;
                10'd817: o_data <= 32'h00009049;
                10'd818: o_data <= 32'h0000913A;
                10'd819: o_data <= 32'h00F08049;
                10'd820: o_data <= 32'h0000904D;
                10'd821: o_data <= 32'h0000912E;
                10'd822: o_data <= 32'h00F0804D;
                10'd823: o_data <= 32'h0000913A;
                10'd824: o_data <= 32'h00F0904B;
                10'd825: o_data <= 32'h0000912E;
                10'd826: o_data <= 32'h00F0804B;
                10'd827: o_data <= 32'h00009049;
                10'd828: o_data <= 32'h0000913A;
                10'd829: o_data <= 32'h00F08049;
                10'd830: o_data <= 32'h00009048;
                10'd831: o_data <= 32'h0000912D;
                10'd832: o_data <= 32'h00F08048;
                10'd833: o_data <= 32'h00009139;
                10'd834: o_data <= 32'h00F08139;
                10'd835: o_data <= 32'h0000912D;
                10'd836: o_data <= 32'h00F09049;
                10'd837: o_data <= 32'h00009139;
                10'd838: o_data <= 32'h00F08049;
                10'd839: o_data <= 32'h0000904B;
                10'd840: o_data <= 32'h00009129;
                10'd841: o_data <= 32'h00F0804B;
                10'd842: o_data <= 32'h00009135;
                10'd843: o_data <= 32'h00F0904D;
                10'd844: o_data <= 32'h00009129;
                10'd845: o_data <= 32'h00F0804D;
                10'd846: o_data <= 32'h00009135;
                10'd847: o_data <= 32'h00F09049;
                10'd848: o_data <= 32'h0000912E;
                10'd849: o_data <= 32'h00F08049;
                10'd850: o_data <= 32'h0000913A;
                10'd851: o_data <= 32'h00F09046;
                10'd852: o_data <= 32'h0000912E;
                10'd853: o_data <= 32'h00F08046;
                10'd854: o_data <= 32'h0000913A;
                10'd855: o_data <= 32'h00F09046;
                10'd856: o_data <= 32'h0000912E;
                10'd857: o_data <= 32'h00F08046;
                10'd858: o_data <= 32'h0000913A;
                10'd859: o_data <= 32'h00F0813A;
                10'd860: o_data <= 32'h00009130;
                10'd861: o_data <= 32'h00F08130;
                10'd862: o_data <= 32'h00009131;
                10'd863: o_data <= 32'h00F08131;
                10'd864: o_data <= 32'h00009133;
                10'd865: o_data <= 32'h00F0904B;
                10'd866: o_data <= 32'h00009127;
                10'd867: o_data <= 32'h00F0804B;
                10'd868: o_data <= 32'h00008127;
                10'd869: o_data <= 32'h00F0904E;
                10'd870: o_data <= 32'h00009127;
                10'd871: o_data <= 32'h00F0804E;
                10'd872: o_data <= 32'h00009052;
                10'd873: o_data <= 32'h00008127;
                10'd874: o_data <= 32'h00F08052;
                10'd875: o_data <= 32'h00009127;
                10'd876: o_data <= 32'h00788127;
                10'd877: o_data <= 32'h00009127;
                10'd878: o_data <= 32'h00789050;
                10'd879: o_data <= 32'h0000912E;
                10'd880: o_data <= 32'h00F08050;
                10'd881: o_data <= 32'h0000904E;
                10'd882: o_data <= 32'h0000912C;
                10'd883: o_data <= 32'h00F0804E;
                10'd884: o_data <= 32'h0000904D;
                10'd885: o_data <= 32'h00009125;
                10'd886: o_data <= 32'h00F0804D;
                10'd887: o_data <= 32'h00009131;
                10'd888: o_data <= 32'h00F08131;
                10'd889: o_data <= 32'h00009125;
                10'd890: o_data <= 32'h00F09049;
                10'd891: o_data <= 32'h00009131;
                10'd892: o_data <= 32'h00F08049;
                10'd893: o_data <= 32'h0000904D;
                10'd894: o_data <= 32'h00009125;
                10'd895: o_data <= 32'h00F0804D;
                10'd896: o_data <= 32'h0000904E;
                10'd897: o_data <= 32'h0000912C;
                10'd898: o_data <= 32'h0078804E;
                10'd899: o_data <= 32'h0000904D;
                10'd900: o_data <= 32'h0078804D;
                10'd901: o_data <= 32'h0000904B;
                10'd902: o_data <= 32'h00009125;
                10'd903: o_data <= 32'h00F0804B;
                10'd904: o_data <= 32'h00009049;
                10'd905: o_data <= 32'h0000912C;
                10'd906: o_data <= 32'h00F08049;
                10'd907: o_data <= 32'h00009048;
                10'd908: o_data <= 32'h0000812C;
                10'd909: o_data <= 32'h00F08048;
                10'd910: o_data <= 32'h01E09049;
                10'd911: o_data <= 32'h00F08049;
                10'd912: o_data <= 32'h0000904B;
                10'd913: o_data <= 32'h00F0804B;
                10'd914: o_data <= 32'h00009045;
                10'd915: o_data <= 32'h00F08045;
                10'd916: o_data <= 32'h0000904D;
                10'd917: o_data <= 32'h00F0804D;
                10'd918: o_data <= 32'h00009045;
                10'd919: o_data <= 32'h00F08045;
                10'd920: o_data <= 32'h00009049;
                10'd921: o_data <= 32'h00F08049;
                10'd922: o_data <= 32'h00F09046;
                10'd923: o_data <= 32'h00F08046;
                10'd924: o_data <= 32'h00F09046;
                10'd925: o_data <= 32'h03C08046;
                10'd926: o_data <= 32'h0000FF2F;
                
                default: o_data <= 32'h0000FF2F;
            endcase
        end
    end

endmodule
